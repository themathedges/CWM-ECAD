//////////////////////////////////////////////////////////////////////////////////
// Test bench for Exercise #5 - Traffic Lights
// Student Name:
// Date: 
//
// Description: A testbench module to test Ex5 - Traffic Lights
// You need to write the whole file
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ns/100ps

module testbench();

parameter clk_period = 10;

reg clk, err;
reg [2:0] prev;
wire [2:0] state;
assign red = state[2];
assign amber = state[1];
assign green = state[0];

initial begin
	clk = 0;
	forever
		#(clk_period/2)clk = ~clk; 		// delay of half a cycle, clk = bitwise not clk 
	end

initial begin	   
	prev = state;
	err = 0;					// prev will hopefully store the previous value of state, in which [111] represents [RAG]
	#clk_period

	forever begin
		#(10*clk_period) 			
		if ((state == 3'b110) && (prev != 3'b100))
		$display("TEST FAILED");
		err = 1;

		if ((state == 3'b001) && (prev != 3'b110))
		$display("TEST FAILED");
		err = 1;

		if ((state == 3'b010) && (prev != 3'b001))
		$display("TEST FAILED");
		err = 1;

		if ((state == 3'b100) && (prev != 3'b010)) //I think I could add a default?
		$display("TEST FAILED");
		err = 1;

		end
end

initial begin
	#(10*clk_period)
	if (err == 0)
	$display("TEST PASSED");				
	$finish;
	end 

traffic traffic(.clk(clk), .red(red), .amber(amber), .green(green)); 		

endmodule 
